entity sm_add_test is
port(
  clk :in std_logic;
  btn : in std_logic_vector (1 downto 0);
  sw : in std_logic_vector (7 downto 0);
  an : out std_logic_vector (3 downto 0);
  sseg : out std_logic_vector (7 downto 0)
);
end sm_add_test;
  
architecture arch_sm of sm_add_test is
signal sum, mout, oct : std_logic_vector (3 downto 0);
signal led3, led2, led1, led0 : std_logic_vector (7 downto 0);
begin
  sm_adder_unit : entity work.sign_mag_add
  generic map(N => 4)
  port map(
    a => sw (3 downto 0),
    b => sw (7 downto 4),
    sum => sum
  );
  with btn select
    mout <= sw (3 downto 0) when "00",
    sw (7 downto 4) when "01",
    sum when others;
  oct <= '0' & mout(2 downto 0);
  sseg_unit : entity work.hex_to_seg
  port map (
    segsig => oct, dp => '1', code_hex => led0);
    led1 <= "10111111" when mout(3) ='1' else "11111111";
    led2 <= "11111111";
    led3 <= "11111111");
  disp_unit:entity work.disp_mux
  port map(
    clk => clk, reset =>'0',
    in0 => led0, in1 => led1, in2 => led2, in3 => led3,
    an => an, sseg => sseg);
end arch_sm;
